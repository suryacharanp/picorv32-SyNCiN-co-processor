module multiplier_bf16(
        input_a,
        input_b,
        mult_input_STB,
        mult_BUSY,
        clk,
        rst,
        output_mult,
        mult_output_STB,
        output_module_BUSY
		);

  input     clk;
  input     rst;

  input     [15:0] input_a;
  input     [15:0] input_b;
  
  input     mult_input_STB;
  output    mult_BUSY;

  output    [15:0] output_mult;
  output    mult_output_STB;
  input     output_module_BUSY;

  //Intermediate registers
  reg       mult_output_STB_reg;
  reg       [15:0] output_mult_reg;
  reg       mult_BUSY_reg;

  reg       [3:0] mult_state;
  parameter get_a_and_b   = 4'd0,
            unpack        = 4'd1,
            special_cases = 4'd2,
            normalise_a   = 4'd3,
            normalise_b   = 4'd4,
            multiply_0    = 4'd5,
            multiply_1    = 4'd6,
            normalise_1   = 4'd7,
            normalise_2   = 4'd8,
            round         = 4'd9,
            pack          = 4'd10,
            put_z         = 4'd11;

  reg       [15:0] a, b, z;
  reg       [7:0] a_m, b_m, z_m;
  reg       [9:0] a_e, b_e, z_e;
  reg       a_s, b_s, z_s;
  reg       guard, round_bit, sticky;
  reg       [49:0] product;

  always @(posedge clk)
  begin

    case(mult_state)

	  
	  get_a_and_b: //Initial state wait for valid inputs and make BUSY = 0 because it has finished previous operation 
      begin
        mult_BUSY_reg <= 0;
        if (!(mult_BUSY_reg) && mult_input_STB) begin  //Once it gets valid input take that input and start processing.
          a <= {input_a};
		  b <= {input_b};
          mult_BUSY_reg <= 1; //Turn the BUSY signal on, BUSY = 1 because now it will be busy processing latched inputs and can no more take inputs even if it is valid. 
          mult_state <= unpack;
        end
      end

      unpack:
      begin
        a_m <= a[6 : 0];
        b_m <= b[6 : 0];
        a_e <= a[14 : 7] - 127;
        b_e <= b[14 : 7] - 127;
        a_s <= a[15];
        b_s <= b[15];
        mult_state <= special_cases;
      end

      special_cases:
      begin
        //if a is NaN or b is NaN return NaN 
        if ((a_e == 128 && a_m != 0) || (b_e == 128 && b_m != 0)) begin
          z[15] <= 1;
          z[14:7] <= 255;
          z[6] <= 1;
          z[5:0] <= 0;
          mult_state <= put_z;
        //if a is inf return inf
        end else if (a_e == 128) begin
          z[15] <= a_s ^ b_s;
          z[14:7] <= 255;
          z[6:0] <= 0;
          //if b is zero return NaN
          if (($signed(b_e) == -127) && (b_m == 0)) begin
            z[15] <= 1;
            z[14:7] <= 255;
            z[6] <= 1;
            z[5:0] <= 0;
          end
          mult_state <= put_z;
        //if b is inf return inf
        end else if (b_e == 128) begin
          z[15] <= a_s ^ b_s;
          z[14:7] <= 255;
          z[6:0] <= 0;
          //if a is zero return NaN
          if (($signed(a_e) == -127) && (a_m == 0)) begin
            z[15] <= 1;
            z[14:7] <= 255;
            z[6] <= 1;
            z[5:0] <= 0;
          end
          mult_state <= put_z;
        //if a is zero return zero
        end else if (($signed(a_e) == -127) && (a_m == 0)) begin
          z[15] <= a_s ^ b_s;
          z[14:7] <= 0;
          z[6:0] <= 0;
          mult_state <= put_z;
        //if b is zero return zero
        end else if (($signed(b_e) == -127) && (b_m == 0)) begin
          z[15] <= a_s ^ b_s;
          z[14:7] <= 0;
          z[6:0] <= 0;
          mult_state <= put_z;
        end else begin
          //Denormalised Number
          if ($signed(a_e) == -127) begin
            a_e <= -126;
          end else begin
            a_m[7] <= 1;
          end
          //Denormalised Number
          if ($signed(b_e) == -127) begin
            b_e <= -126;
          end else begin
            b_m[7] <= 1;
          end
          mult_state <= normalise_a;
        end
      end

      normalise_a:
      begin
        if (a_m[7]) begin
          mult_state <= normalise_b;
        end else begin
          a_m <= a_m << 1;
          a_e <= a_e - 1;
        end
      end

      normalise_b:
      begin
        if (b_m[7]) begin
          mult_state <= multiply_0;
        end else begin
          b_m <= b_m << 1;
          b_e <= b_e - 1;
        end
      end

      multiply_0:
      begin
        z_s <= a_s ^ b_s;
        z_e <= a_e + b_e + 1;
        product <= a_m * b_m * 4;
        mult_state <= multiply_1;
      end

      multiply_1:
      begin
        z_m <= product[49:26];
        guard <= product[25];
        round_bit <= product[24];
        sticky <= (product[23:0] != 0);
        mult_state <= normalise_1;
      end

      normalise_1:
      begin
        if (z_m[7] == 0) begin
          z_e <= z_e - 1;
          z_m <= z_m << 1;
          z_m[0] <= guard;
          guard <= round_bit;
          round_bit <= 0;
        end else begin
          mult_state <= normalise_2;
        end
      end

      normalise_2:
      begin
        if ($signed(z_e) < -126) begin
          z_e <= z_e + 1;
          z_m <= z_m >> 1;
          guard <= z_m[0];
          round_bit <= guard;
          sticky <= sticky | round_bit;
        end else begin
          mult_state <= round;
        end
      end

      round:
      begin
        if (guard && (round_bit | sticky | z_m[0])) begin
          z_m <= z_m + 1;
          if (z_m == 8'hff) begin
            z_e <=z_e + 1;
          end
        end
        mult_state <= pack;
      end

      pack:
      begin
        z[6 : 0] <= z_m[6:0];
        z[14 : 7] <= z_e[7:0] + 127;
        z[15] <= z_s;
        if ($signed(z_e) == -126 && z_m[7] == 0) begin
          z[14 : 7] <= 0;
        end
        //if overflow occurs, return inf
        if ($signed(z_e) > 127) begin
          z[6 : 0] <= 0;
          z[14 : 7] <= 255;
          z[15] <= z_s;
        end
        mult_state <= put_z;
      end
	  
	  put_z: //Final state valid output is ready , make the output STB/VALID = 1, put valid output.
      begin
        mult_output_STB_reg <= 1;
        output_mult_reg <= z;
        if (mult_output_STB_reg && !(output_module_BUSY)) begin //Once output module is no more BUSY it lowers it's busy signal and output is then taken by next module.
          mult_output_STB_reg <= 0; //Output is no more valid.
          mult_state <= get_a_and_b; //Go back to initial state.
        end
      end

    endcase

	
	 if (rst == 1) begin //At Active high reset, module is no more BUSY, go to initial state and wait for valid inputs. Input is don't care and output is don't care , so output VALID/STB = 0.
      mult_state <= get_a_and_b;
      mult_BUSY_reg <= 0; 
      mult_output_STB_reg <= 0;
    end

  end
  
  
   `ifdef SYNTHESIS_OFF //Purely combinational logic for debugging purpose, based on hexadecimal encoded states it will show named states in waveform 
   //see this register "statename" in ASCII in dump
  reg [8*13:0] mult_statename;//Highest 13 Number of ASCII letters each 8 bits.
  always@* begin
    case (1'b1)
      (mult_state === get_a_and_b)  : mult_statename = "GET_A_AND_B";
      (mult_state === unpack)       : mult_statename = "UNPACK";
      (mult_state === special_cases): mult_statename = "SPECIAL_CASES";//13 ASCII letters
      (mult_state === normalise_a)  : mult_statename = "NORMALISE_A";
      (mult_state === normalise_b)  : mult_statename = "NORMALISE_B";
      (mult_state === multiply_0)   : mult_statename = "MULTIPLY_0";
      (mult_state === multiply_1)   : mult_statename = "MULTIPLY_1";
      (mult_state === normalise_1)  : mult_statename = "NORMALIZE_1";
      (mult_state === normalise_2)  : mult_statename = "NORMALIZE_2";
      (mult_state === round)        : mult_statename = "ROUND";
      (mult_state === pack)         : mult_statename = "PACK";
      (mult_state === put_z)        : mult_statename = "PUT_Z";
    endcase
  end//always
  `endif
  
  

  //Continuous assignments
  
  assign mult_BUSY = mult_BUSY_reg;
  assign mult_output_STB = mult_output_STB_reg;
  assign output_mult = output_mult_reg[31:16];

endmodule : multiplier